This is a test for hl setting
