lcls
lmc
lmhelp
int val0
int val1
