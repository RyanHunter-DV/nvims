lcls
lmc
lmhelp
int val0
int val1
cld
function void build_phase (uvm_phase phase);
endfunction
